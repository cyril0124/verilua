module Design (
    input wire clock,
    input wire reset,
    input reg [15:0]  value16,
    input reg [31:0]  value32,
    input reg [63:0]  value64,
    input reg [127:0] value128
);  

endmodule