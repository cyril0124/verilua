module Design (
    input wire clock,
    input wire reset,
    input wire [15:0]  value16,
    input wire [31:0]  value32,
    input wire [63:0]  value64,
    input wire [127:0] value128
);  

endmodule